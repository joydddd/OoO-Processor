`timescale 1ns/100ps
`ifndef __PIPELINE_TEST_SV__
`define __PIPELINE_TEST_SV__

`define TEST_MODE 
`define DIS_DEBUG
`define CACHE_MODE
`define CACHE_SIM // TODO: comment this line to use real cache instead of simulation

/* import freelist simulator */
import "DPI-C" function void fl_init();
import "DPI-C" function int fl_new_pr_valid();
import "DPI-C" function int fl_new_pr2(int new_pr_en);
import "DPI-C" function int fl_new_pr1(int new_pr_en);
import "DPI-C" function int fl_new_pr0(int new_pr_en);
import "DPI-C" function int fl_pop(int new_pr_en);

/* import map table simulator */ 
import "DPI-C" function void mt_init();
import "DPI-C" function int mt_look_up(int i);
import "DPI-C" function int mt_look_up_ready(int i);
import "DPI-C" function void mt_map(int ar, int pr);

/* import print pipeline */
import "DPI-C" function void print_header(string str);
import "DPI-C" function void print_num(int num);
import "DPI-C" function void print_stage(string div, int inst, int npc, int valid_inst);

/* import print rs */ 
import "DPI-C" function void print_select(int index,  int valid, int inst,  int npc, int fu_select, int op_select);

/* import simulate cache & memory */
import "DPI-C" function void mem_init();
import "DPI-C" function void mem_write(int addr, int data, int byte3, byte2, byte1, byte0);
import "DPI-C" function int mem_read(int addr);
import "DPI-C" function void mem_print();

module testbench;
logic clock, reset;

`ifdef TEST_MODE
// IF to Dispatch 


// ID stage output
IF_ID_PACKET [2:0]         dis_in_display;
ROB_ENTRY_PACKET [2:0]     dis_rob_packet_display;
logic [2:0]                dis_stall_display;

// RS
RS_IN_PACKET [2:0]         dis_rs_packet_display;
RS_IN_PACKET [`RSW-1:0]    rs_entries_display;
RS_S_PACKET [2:0]          rs_out_display;
logic [2:0]                rs_stall_display;

// Maptable
logic [31:0][`PR-1:0] map_array_display;
logic [31:0] ready_array_display;
logic [31:0][`PR-1:0] archi_map_display;

// IS
RS_S_PACKET [2:0]          is_in_display;
FU_FIFO_PACKET             fu_fifo_stall_display;
ISSUE_FU_PACKET [`IS_FIFO_DEPTH-1:0] alu_fifo_display;
ISSUE_FU_PACKET [`IS_FIFO_DEPTH-1:0] mult_fifo_display;
ISSUE_FU_PACKET [`IS_FIFO_DEPTH-1:0] br_fifo_display;
ISSUE_FU_PACKET [`IS_FIFO_DEPTH-1:0] ls_fifo_display;


// FU 
ISSUE_FU_PACKET [2**`FU-1:0] fu_in_display;
FU_STATE_PACKET            fu_ready_display;
FU_STATE_PACKET            fu_finish_display;
FU_COMPLETE_PACKET [2**`FU-1:0]   fu_packet_out_display;

// SQ
SQ_ENTRY_PACKET [0:2**`LSQ-1]  sq_display;
logic [`LSQ-1:0]               head_dis;
logic [`LSQ-1:0]               tail_dis;
logic [`LSQ:0]                 filled_num_dis;
SQ_ENTRY_PACKET [2**`LSQ-1:0]  older_stores;
logic [2**`LSQ-1:0]            older_stores_valid;
LOAD_SQ_PACKET [1:0]           load_sq_pckt_display;

// Complete
CDB_T_PACKET               cdb_t_display;
FU_COMPLETE_PACKET [2:0]    complete_pckt_in_display;
logic [2**`FU-1:0]          complete_stall_display;

//ROB
	ROB_ENTRY_PACKET [`ROBW-1:0]    rob_entries_display;
    logic       [`ROB-1:0]          head_display;
    logic       [`ROB-1:0]          tail_display;
    logic       [2:0]               rob_stall_display;

// PR
    logic [2**`PR-1:0][`XLEN-1:0] pr_display;

// Archi Map Table
    logic [2:0][`PR-1:0]       map_ar_pr;
    logic [2:0][4:0]           map_ar;

    logic [31:0][`PR-1:0]            fl_array_display;
    logic [4:0]                      fl_head_display;
    logic [4:0]                      fl_tail_display;
    logic                            fl_empty_display;

`endif

`ifdef DIS_DEBUG
IF_ID_PACKET [2:0]          if_d_packet_debug;
logic [2:0]                 dis_new_pr_en_out;
/* free list simulation */
logic [2:0]                 free_pr_valid_debug;
logic [2:0][`PR-1:0]        free_pr_debug;

/* maptable simulation */
/*
logic [2:0] [4:0]           maptable_lookup_reg1_ar_out;
logic [2:0] [4:0]           maptable_lookup_reg2_ar_out;
logic [2:0] [4:0]           maptable_allocate_ar_out;
logic [2:0] [`PR-1:0]       maptable_allocate_pr_out;
logic [2:0][`PR-1:0]        maptable_old_pr_debug;
logic [2:0][`PR-1:0]        maptable_reg1_pr_debug;
logic [2:0][`PR-1:0]        maptable_reg2_pr_debug;
logic [2:0]                 maptable_reg1_ready_debug;
logic [2:0]                 maptable_reg2_ready_debug;
*/

logic [2:0]                 rob_stall_debug;
FU_STATE_PACKET             fu_ready_debug;
CDB_T_PACKET                cdb_t_debug;
`endif


SQ_ENTRY_PACKET [2:0]          cache_wb_sim;
logic [1:0][`XLEN-1:0]         cache_read_addr_sim;
logic [1:0][`XLEN-1:0]         cache_read_data_sim;
logic [1:0]                    cache_read_start_sim;

logic  [3:0]        Imem2proc_response;
logic [63:0]        Imem2proc_data;
logic  [3:0]        Imem2proc_tag;
logic [`XLEN-1:0]   proc2Imem_addr;
logic [1:0]         proc2Imem_command;

mem memory(
    .clk(clock),                            // Memory clock
    .proc2mem_addr(proc2Imem_addr),         // <- pipeline.proc2mem_addr
    //support for memory model with byte level addressing
    // TODO: change when we have store and load
    .proc2mem_data(64'b0),                  // write data, no need for this test 
`ifndef CACHE_MODE  
    .proc2mem_size(DOUBLE),                 //BYTE, HALF, WORD or DOUBLE, no need for this test
`endif
    // TODO: when we have store and load FU, this signal connection needs to be modified
    .proc2mem_command(proc2Imem_command),   // `BUS_NONE `BUS_LOAD or `BUS_STORE
    
    .mem2proc_response(Imem2proc_response), // 0 = can't accept, other=tag of transaction
    .mem2proc_data(Imem2proc_data),         // data resulting from a load
    .mem2proc_tag(Imem2proc_tag)            // 0 = no value, other=tag of transaction
);

pipeline tbd(
    .clock(clock),
    .reset(reset),
    .mem2proc_response(Imem2proc_response),    // <- mem.mem2proc_response
	.mem2proc_data(Imem2proc_data),            // <- mem.mem2proc_data
	.mem2proc_tag(Imem2proc_tag),              // <- mem.mem2proc_tag
	
	.proc2mem_command(proc2Imem_command),      // -> mem.proc2Imem_command
	.proc2mem_addr(proc2Imem_addr)             // -> mem.proc2Imem_addr
`ifdef TEST_MODE
    // ID
    , .dis_in_display(dis_in_display)
    , .dis_rob_packet_display(dis_rob_packet_display)
    , .dis_stall_display(dis_stall_display)
    // RS
    , .dis_rs_packet_display(dis_rs_packet_display)
    , .rs_entries_display(rs_entries_display)
    , .rs_out_display(rs_out_display)
    , .rs_stall_display(rs_stall_display)
    // Maptable
    , .map_array_disp(map_array_display)
    , .ready_array_disp(ready_array_display)
    , .archi_map_display(archi_map_display)
    // IS
    , .is_in_display(is_in_display)
    , .fu_fifo_stall_display(fu_fifo_stall_display)
    , .alu_fifo_display(alu_fifo_display)
    , .mult_fifo_display(mult_fifo_display)
    , .br_fifo_display(br_fifo_display)
    , .ls_fifo_display(ls_fifo_display)
    // FU
    , .fu_in_display(fu_in_display)
    , .fu_ready_display(fu_ready_display)
    , .fu_finish_display(fu_finish_display)
    , .fu_packet_out_display(fu_packet_out_display)
    // SQ
    , .sq_display(sq_display)
    , .head_dis(head_dis)
    , .tail_dis(tail_dis)
    , .filled_num_dis(filled_num_dis)
    , .older_stores(older_stores)
    , .older_stores_valid(older_stores_valid)
    , .load_sq_pckt_display(load_sq_pckt_display)
    // Complete
    , .cdb_t_display(cdb_t_display)
    , .wb_value_display(wb_value_display)
    , .complete_pckt_in_display(complete_pckt_in_display)
    , .complete_stall_display(complete_stall_display)
    // ROB
    , .rob_entries_display(rob_entries_display)
    , .head_display(head_display)
    , .tail_display(tail_display)
    , .rob_stall_display(rob_stall_display)
    // Freelist
    , .fl_array_display(fl_array_display)
    , .fl_head_display(fl_head_display)
    , .fl_tail_display(fl_tail_display)
    , .fl_empty_display(fl_empty_display)
    // PR
    , .pr_display(pr_display)
    // Archi Map Table
    , .map_ar_pr_disp(map_ar_pr)
    , .map_ar_disp(map_ar)
`endif // TEST_MODE

`ifdef DIS_DEBUG
    , .if_d_packet_debug(if_d_packet_debug)
    , .dis_new_pr_en_out(dis_new_pr_en_out)
    /* free list simulation */
    // , .free_pr_valid_debug(free_pr_valid_debug)
    // , .free_pr_debug(free_pr_debug)
    /* maptable simulation */
    /*
    , .maptable_lookup_reg1_ar_out(maptable_lookup_reg1_ar_out)
    , .maptable_lookup_reg2_ar_out(maptable_lookup_reg2_ar_out)
    , .maptable_allocate_ar_out(maptable_allocate_ar_out)
    , .maptable_allocate_pr_out(maptable_allocate_pr_out)
    , .maptable_old_pr_debug(maptable_old_pr_debug)
    , .maptable_reg1_pr_debug(maptable_reg1_pr_debug)
    , .maptable_reg2_pr_debug(maptable_reg2_pr_debug)
    , .maptable_reg1_ready_debug(maptable_reg1_ready_debug)
    , .maptable_reg2_ready_debug(maptable_reg2_ready_debug)
    */

    // , .rob_stall_debug(rob_stall_debug)
    // , .fu_ready_debug(fu_ready_debug)
    // , .cdb_t_debug(cdb_t_debug)
`endif
`ifdef CACHE_SIM
    , .cache_wb_sim(cache_wb_sim)
    , .cache_read_addr_sim(cache_read_addr_sim)
    , .cache_read_data_sim(cache_read_data_sim)
    , .cache_read_start_sim(cache_read_start_sim)
`endif
);

/* clock */
always begin
	#(`VERILOG_CLOCK_PERIOD/2.0);
	clock = ~clock;
end

////////////////////////////////////////////////////////////
/////////////       SIMULATORS
///////////////////////////////////////////////////////////

int cycle_count; 
always @(posedge clock) begin
    cycle_count++;
end

`ifdef CACHE_SIM
always @(posedge clock) begin
    if (reset) begin
        mem_init();
    end
end

always @(posedge clock) begin
    if (!reset) begin
        mem_write(cache_wb_sim[0].addr, cache_wb_sim[0].data, cache_wb_sim[0].usebytes[3], cache_wb_sim[0].usebytes[2], cache_wb_sim[0].usebytes[1], cache_wb_sim[0].usebytes[0]);
        mem_write(cache_wb_sim[1].addr, cache_wb_sim[1].data, cache_wb_sim[1].usebytes[3], cache_wb_sim[1].usebytes[2], cache_wb_sim[1].usebytes[1], cache_wb_sim[1].usebytes[0]);
        mem_write(cache_wb_sim[2].addr, cache_wb_sim[2].data, cache_wb_sim[2].usebytes[3], cache_wb_sim[2].usebytes[2], cache_wb_sim[2].usebytes[1], cache_wb_sim[2].usebytes[0]);
    end
end

always @(cache_read_addr_sim, cache_read_start_sim) begin
    if (cache_read_start_sim[0]) cache_read_data_sim[0] = mem_read(cache_read_addr_sim[0]);
    if (cache_read_start_sim[1]) cache_read_data_sim[1] = mem_read(cache_read_addr_sim[1]);
end

`endif
// /* free list simulator */
// always @(posedge clock) begin
//     if (reset) begin
//         fl_init();
//     end else begin
//         fl_pop(dis_new_pr_en_out);
//     end
// end
// always @(dis_new_pr_en_out, clock) begin
//     `SD;
//     if (!reset) begin
//         free_pr_valid_debug = fl_new_pr_valid();
//         free_pr_debug[2] = fl_new_pr2(dis_new_pr_en_out);
//         free_pr_debug[1] = fl_new_pr1(dis_new_pr_en_out);
//         free_pr_debug[0] = fl_new_pr0(dis_new_pr_en_out);
//     end
// end

/* map table simulator */
/*
always @(posedge clock) begin
    if (reset) begin
        mt_init();
    end else begin
        for(int i=0; i<3; i++) begin
            mt_map(maptable_allocate_ar_out[i], maptable_allocate_pr_out[i]); 
        end
    end
end
always @(maptable_allocate_ar_out) begin
    maptable_old_pr_debug[2] = mt_look_up(maptable_allocate_ar_out[2]);
    maptable_old_pr_debug[1] = mt_look_up(maptable_allocate_ar_out[1]);
    maptable_old_pr_debug[0] = mt_look_up(maptable_allocate_ar_out[0]);
end
always @(maptable_lookup_reg1_ar_out) begin
    for(int i=0; i<3; i++) begin
        maptable_reg1_pr_debug[i] = mt_look_up(maptable_lookup_reg1_ar_out[i]);
        maptable_reg1_ready_debug[i] = mt_look_up_ready(maptable_lookup_reg1_ar_out[i]);
    end
end
always @(maptable_lookup_reg2_ar_out) begin
    for(int i=0; i<3; i++) begin
        maptable_reg2_pr_debug[i] = mt_look_up(maptable_lookup_reg2_ar_out[i]);
        maptable_reg2_ready_debug[i] = mt_look_up_ready(maptable_lookup_reg2_ar_out[i]);
    end
end

*/

//////////////////////////////////////////////////////////////
//////////////                  DISPLAY
/////////////////////////////////////////////////////////////
always @(negedge clock) begin
    if (!reset)  begin
        #1;
        print_retire_wb();
        // $display();
        // $display("~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~");
        // $display();
        
        if (cycle_count >= 500 && cycle_count <= 520) print_pipeline;
        if (cycle_count >= 500 && cycle_count <= 520) print_alu;
        // show_fu_stat;
        // print_is_fifo;
        // show_sq;
        // show_sq_age;
        // show_cdb;
        // show_rs_in;
        
        // show_complete;
        if (cycle_count >= 500 && cycle_count <= 520) show_rs_table;
        if (cycle_count >= 510 && cycle_count <= 520) show_rob_table;
        // show_rob_in;
        // show_rs_out;
        // show_freelist_table;
        // show_mpt_entry;
    end
end


task show_rs_in;
    begin
        $display("=====   RS_IN Packet   =====");
        $display("| WAY |     inst    | fu_sel | op_sel  |");
        for (int i=2; i >= 0 ; i--) begin
            print_select(i, dis_rs_packet_display[i].valid, dis_rs_packet_display[i].inst, dis_rs_packet_display[i].PC, dis_rs_packet_display[i].fu_sel, dis_rs_packet_display[i].op_sel);
        end
        $display("| WAY | dest_pr | reg1_pr | reg1_ready | reg2_pr | reg2_ready |");
        for (int i=2; i>=0; i--) begin
            $display("|  %1d  |      %2d |      %2d |          %b |     %2d  |          %b |",
                i, dis_rs_packet_display[i].dest_pr, dis_rs_packet_display[i].reg1_pr, dis_rs_packet_display[i].reg1_ready, dis_rs_packet_display[i].reg2_pr, dis_rs_packet_display[i].reg2_ready
            );
        end
    end
endtask

task show_rs_out;
    begin
        $display("=====   RS_S Packet   =====");
        $display("| WAY |     inst    | fu_sel | op_sel  |");
        for (int i=2; i>=0; i--) begin
            print_select(i, rs_out_display[i].valid, rs_out_display[i].inst, rs_out_display[i].PC, rs_out_display[i].fu_sel, rs_out_display[i].op_sel);
        end
        $display("| WAY | valid |  PC  | dest_pr | reg1_pr | reg2_pr |       inst | halt |");
        for (int i=2; i>=0; i--) begin
            $display("|  %1d  |     %b | %4h |      %2d |      %2d |     %2d  |",
                i, rs_out_display[i].valid, rs_out_display[i].PC, rs_out_display[i].dest_pr, rs_out_display[i].reg1_pr, rs_out_display[i].reg2_pr, rs_out_display[i].inst, rs_out_display[i].halt
            );
        end
    end
endtask

task show_rs_table;
    for(int i=2**`RS-1; i>=0; i--) begin  // For RS entry, it allocates from 15-0
        print_stage("*", rs_entries_display[i].inst, rs_entries_display[i].PC[31:0], rs_entries_display[i].valid);
        $display("dest_pr:%d reg1_pr:%d reg1_ready: %b reg2_pr:%d reg2_ready %b rob_entry:%d", rs_entries_display[i].dest_pr, rs_entries_display[i].reg1_pr, rs_entries_display[i].reg1_ready, rs_entries_display[i].reg2_pr, rs_entries_display[i].reg2_ready, rs_entries_display[i].rob_entry);
    end
    $display("structual_stall:%b", rs_stall_display);
endtask; // show_rs_table


task show_fu_stat;
    $display("fu ready: %8b", fu_ready_display);
    $display("fu finish: %8b", fu_finish_display);
    $display("| valid | halt | take_branch | target_pc | dest_pr | dest_value | rob_entry |");
    for(int i=0; i<2**`FU; i++) begin
        $display("| %1d | %1d | %1d | %4h | %2d | %d | %2d |", 
                fu_packet_out_display[i].valid, fu_packet_out_display[i].halt, fu_packet_out_display[i].if_take_branch,
                fu_packet_out_display[i].target_pc, fu_packet_out_display[i].dest_pr, fu_packet_out_display[i].dest_value,
                fu_packet_out_display[i].rob_entry);
    end
endtask; 

task show_sq;
    $display("HEAD: %d, Tail: %d, Filled num: %d", head_dis, tail_dis, filled_num_dis);
    $display(" |ready|   addr   |usebytes|   data   |");
    for(int i=0; i<2**`LSQ; i++) begin
        $display("%1d|  %d  | %8h |  %4b  | %8h |", i, sq_display[i].ready, sq_display[i].addr, sq_display[i].usebytes, sq_display[i].data);
    end
endtask

task show_sq_age;
    $display("##### older stores, tail_pos at %d", load_sq_pckt_display[0].tail_pos);
    $display(" |valid|ready|   addr   |usebytes|   data   |");
    for(int i=0; i<2**`LSQ; i++) begin
        $display("%1d|  %d  |  %d  | %8h |  %4b  | %8h |", i, older_stores_valid[i], older_stores[i].ready, older_stores[i].addr, older_stores[i].usebytes, older_stores[i].data);
    end
endtask


task show_complete;
    $display("fu ready: %8b", fu_ready_display);
    $display("complete stall: %8b", complete_stall_display);
    $display("======== Completing =============");
    $display("| valid | halt | take_branch | target_pc | dest_pr | dest_value | rob_entry |");
    for(int i=0; i<3; i++) begin
        $display("| %1d | %1d | %1d | %4h | %2d | %d | %2d |", 
                complete_pckt_in_display[i].valid, complete_pckt_in_display[i].halt, complete_pckt_in_display[i].if_take_branch,
                complete_pckt_in_display[i].target_pc, complete_pckt_in_display[i].dest_pr, complete_pckt_in_display[i].dest_value,
                complete_pckt_in_display[i].rob_entry);
    end
endtask; 

task show_cdb;
    $display("CDB: %d  %d  %d", cdb_t_display.t0, cdb_t_display.t1, cdb_t_display.t2);
endtask;

task show_rob_in;
    $display("|ROB|valid| Tnew | Told | Reg  |Completed|");
    for(int i=2; i>=0; i--) begin
        $display("| %1d |  %1d  |  %2d  |  %2d  |  %2d  |    %1d    |", i, dis_rob_packet_display[i].valid, dis_rob_packet_display[i].Tnew, dis_rob_packet_display[i].Told, dis_rob_packet_display[i].arch_reg, dis_rob_packet_display[i].completed);
    end
endtask

task show_rob_table;
    for(int i=2**`ROB-1; i>=0; i--) begin  
        $display("%d| valid: %d  Tnew: %d  Told: %d  arch_reg: %d  completed: %b  precise_state: %b  target_pc: %3d is_store: %b", i, rob_entries_display[i].valid, rob_entries_display[i].Tnew, rob_entries_display[i].Told, rob_entries_display[i].arch_reg, rob_entries_display[i].completed, rob_entries_display[i].precise_state_need, rob_entries_display[i].target_pc, rob_entries_display[i].is_store);
    end
    $display("head:%d tail:%d", head_display, tail_display);
    $display("structual_stall:%b", rob_stall_display);
endtask; // show_rs_table


task print_pipeline;
    $display(" ============ Cycle %d ==============", cycle_count);
    print_header("\n |     IF      |     DIS     |     IS      |\n");
    for(int i=2; i>=0; i--) begin
        print_num(i);
        `ifdef DIS_DEBUG
        /* IF debug */
        print_stage("|", if_d_packet_debug[i].inst, if_d_packet_debug[i].PC, if_d_packet_debug[i].valid);
        `endif
        /* DIS */
        print_stage("|", dis_in_display[i].inst, dis_in_display[i].PC, dis_in_display[i].valid);
        // /* dispatch to rs */
        // print_stage("|", dis_rs_packet_display[i].inst, dis_rs_packet_display[i].PC, dis_rs_packet_display[i].valid);
        /* IS */
        print_stage("|", is_in_display[i].inst, is_in_display[i].PC, is_in_display[i].valid);
        print_header("|\n");
    end
    for(int i=2; i>=0; i--) begin
        `ifdef DIS_DEBUG
        /* IF debug */
        $display("%h", if_d_packet_debug[i].inst);
        `endif
    end
endtask

task print_final;
    $display("+++++++++++++++++++++ Result ++++++++++++++++++++++");
    $display("Arch Map Table");
    $display("|  AR  |  PR  |");
    for(int i=0; i<32; i++)begin
        $display("|  %2d  |  %2d  |", i, archi_map_display[i]);
    end
    $display("Physical Register");
    $display("|  PR  |  value  |");
    for(int i=0; i<64; i++)begin
        $display("|  %2d  |  %10d  |", i, pr_display[i]);
    end
    `ifdef CACHE_SIM
    mem_print();
    `endif
endtask

task print_retire_wb;
    for(int i=2; i>=0; i--) begin
        if (map_ar[i] != 0) $display("Cycle: %d: wb r%d = %d", cycle_count, map_ar[i], $signed(pr_display[map_ar_pr[i]]));
    end
endtask
task print_is_fifo;
    $display("IS FIFO stall: %4b", fu_fifo_stall_display);
    print_header("\n|     ALU     |     LS      |    MULT     |   BRANCH    |\n");
    for(int i=0; i<`IS_FIFO_DEPTH; i++) begin
        print_stage("|", alu_fifo_display[i].inst, alu_fifo_display[i].PC, alu_fifo_display[i].valid);
        print_stage("|", ls_fifo_display[i].inst, ls_fifo_display[i].PC, ls_fifo_display[i].valid);
        print_stage("|", mult_fifo_display[i].inst, mult_fifo_display[i].PC, mult_fifo_display[i].valid);
        print_stage("|", br_fifo_display[i].inst, br_fifo_display[i].PC, br_fifo_display[i].valid);
        print_header("|\n");
    end
endtask

task print_alu;
    print_header("\n|    ALU_1    |    ALU_2    |    ALU_3    |     LS_1    |     LS_2    |    MULT_1   |    MULT_2   |    BRANCH   |\n");
    for (int i=0; i<2**`FU; i++) begin
        print_stage("|", fu_in_display[i].inst, fu_in_display[i].PC, fu_in_display[i].valid);
    end
    $display();
endtask

task show_freelist_table;
    for(int i=31; i>=0; i--) begin  // For RS entry, it allocates from 15-0
        $display("Index: %d        PR: %5d", i, fl_array_display[i]);
    end
    $display("head:%d tail:%d empty:%d", fl_head_display, fl_tail_display, fl_empty_display);
endtask; // show_rs_table

task show_mpt_entry;
    begin
        $display("=====   Maptable Entry   =====");
        $display("| AR |   PR   | ready |");
        for (int i = 0; i < 32; i++) begin
            $display("| %2d |   %d   |   %b  |", i, archi_map_display[i], ready_array_display[i]);
        end
        $display(" ");
    end
endtask

//////////////////////////////////////////////////////////
///////////////         SET      
/////////////////////////////////////////////////////////

// task set_if_d_packet;
//     input int i;
//     input INST inst;
//     input [`XLEN-1:0] pc;
//     if_d_packet_debug[i].inst = inst;
//     if_d_packet_debug[i].PC = pc;
//     if_d_packet_debug[i].NPC = pc+4;
//     if_d_packet_debug[i].valid = 1;
// endtask

task set_if_d_packet_invalid;
    input int i;
    if_d_packet_debug[i].valid = 0;
endtask

// int PC; 
initial begin
    $dumpvars;
    clock = 1'b0;
    reset = 1'b1;
    cycle_count = 0;
    // rob_stall_debug = 3'b000;
    // fu_ready_debug = 8'b00011111;
    // cdb_t_debug = {`RS'b0, `RS'b0, `RS'b0};
    // PC = 0;
    @(posedge clock)
    $readmemh("program.mem", memory.unified_memory);
    @(posedge clock)
    #2 reset = 1'b0;
    

    for (int i = 0; i < 750; i++) begin
    @(negedge clock);
    end
    
    #2;
    print_final;
    $display("@@@Pass: test finished");
    $finish;
end

endmodule




`endif // __PIPELINE_TEST_SV__